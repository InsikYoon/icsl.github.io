module PriorityBasedArbiter (


);


end